library verilog;
use verilog.vl_types.all;
entity rxTest_vlg_vec_tst is
end rxTest_vlg_vec_tst;
