library verilog;
use verilog.vl_types.all;
entity uartProject_vlg_vec_tst is
end uartProject_vlg_vec_tst;
