library verilog;
use verilog.vl_types.all;
entity generalTest_vlg_vec_tst is
end generalTest_vlg_vec_tst;
